`ifndef _CPU_SVH_
`define _CPU_SVH_

// シミュレーション設定
`define LOG_PC

`endif // _CPU_SVH_