`ifndef _CPU_SVH_
`define _CPU_SVH_

// シミュレーション設定
`define LOG_PC
`define LOG_IMEM
`define LOG_DECODER
`define LOG_GPR

`endif // _CPU_SVH_